package router_test_pkg;

        import uvm_pkg::*;

        `include "uvm_macros.svh"

        `include "write_xtn.sv"
        `include "wr_agent_config.sv"
        `include "rd_agent_config.sv"
        `include "router_env_config.sv"
        `include "wr_driver.sv"
        `include "wr_monitor.sv"
        `include "wr_sequencer.sv"
        `include "wr_agent.sv"
        `include "wr_agent_top.sv"
        `include "wr_seqs.sv"

        `include "read_xtn.sv"
        `include "rd_monitor.sv"
        `include "rd_sequencer.sv"
        `include "rd_seqs.sv"
        `include "rd_driver.sv"
        `include "rd_agent.sv"
        `include "rd_agent_top.sv"

        `include "router_virtual_sequencer.sv"
        `include "router_virtual_seqs.sv"
        `include "router_scoreboard.sv"

        `include "router_env.sv"


        `include "router_vtest_lib.sv"

endpackage

